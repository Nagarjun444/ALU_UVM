
class alu_monitor extends uvm_monitor;
  `uvm_component_utils(alu_monitor)
  
  virtual alu_interface vif;
   alu_sequence_item item;

  uvm_analysis_port#(alu_sequence_item)monitor_port; // from moniter to scoreboard
   
  
  function new(string name="alu_monitor",uvm_component parent);
     super.new(name,parent);
	 `uvm_info("MONITOR_CLASS","Inside constructor!",UVM_HIGH)
  endfunction
  
  
  //--BUILD PHASE
  
  function void build_phase(uvm_phase phase);
   super.build_phase(phase);
   monitor_port=new("monitor_port",this);                                     // for analysis port we are creating method
   `uvm_info("MONITOR_CLASS","Build phase!",UVM_HIGH)
           
    if(!(uvm_config_db #(virtual alu_interface)::get(this,"*","vif",vif)))
	     begin		   
	     `uvm_error("MONITOR_CLASS","failed to get VIF from calling DBI")
		 end
  endfunction
  
  ///---CONNECT PHASE
  function void connect_phase(uvm_phase phase);
   super.connect_phase(phase);
   `uvm_info("MONITOR_CLASS","Connect phase!",UVM_HIGH)
  endfunction
  
  
  //-----RUN PHASE
  task run_phase(uvm_phase phase);
   begin
    super.run_phase(phase);
	`uvm_info("MONITOR_CLASS","Inside Run phase!",UVM_HIGH)
	
	   //logic
	     forever 
		  begin
		     item = alu_sequence_item::type_id::create("item");
			  wait(!vif.reset);
			   //sample input
			   @(posedge vif.clock);
			       item.a=vif.a;
			       item.b=vif.b;
			       item.op_code=vif.op_code;
				  
				  //sample output
				   @(posedge vif.clock);
				     item.result= vif.result;
					 
					 
					 
					//send item to scoreboard
					monitor_port.write(item);
					
		  end
	end	  
  endtask
endclass


/*

class alu_monitor extends uvm_monitor;
  `uvm_component_utils(alu_monitor)
  
  virtual alu_interface vif;
  alu_sequence_item item;
  
  uvm_analysis_port #(alu_sequence_item) monitor_port;
  
  
  //--------------------------------------------------------
  //Constructor
  //--------------------------------------------------------
  function new(string name = "alu_monitor", uvm_component parent);
    super.new(name, parent);
    `uvm_info("MONITOR_CLASS", "Inside Constructor!", UVM_HIGH)
  endfunction: new
  
  
  //--------------------------------------------------------
  //Build Phase
  //--------------------------------------------------------
  function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    `uvm_info("MONITOR_CLASS", "Build Phase!", UVM_HIGH)
    
    monitor_port = new("monitor_port", this);
    
    if(!(uvm_config_db #(virtual alu_interface)::get(this, "*", "vif", vif))) begin
      `uvm_error("MONITOR_CLASS", "Failed to get VIF from config DB!")
    end
    
  endfunction: build_phase
  
  //--------------------------------------------------------
  //Connect Phase
  //--------------------------------------------------------
  function void connect_phase(uvm_phase phase);
    super.connect_phase(phase);
    `uvm_info("MONITOR_CLASS", "Connect Phase!", UVM_HIGH)
    
  endfunction: connect_phase
  
  
  //--------------------------------------------------------
  //Run Phase
  //--------------------------------------------------------
  task run_phase (uvm_phase phase);
    super.run_phase(phase);
    `uvm_info("MONITOR_CLASS", "Inside Run Phase!", UVM_HIGH)
    
    forever begin
      item = alu_sequence_item::type_id::create("item");
      
      wait(!vif.reset);
      
      //sample inputs
      @(posedge vif.clock);
      item.a = vif.a;
      item.b = vif.b;
      item.op_code = vif.op_code;
      
      //sample output
      @(posedge vif.clock);
      item.result = vif.result;
      
      // send item to scoreboard
      monitor_port.write(item);
    end
        
  endtask: run_phase
  
  
endclass: alu_monitor*/